----------------------------------------------------------------------------------
-- Engineer: 	   Matjaz Mav
-- Create Date:    02/04/2017 
-- Module Name:    canvas - Behavioral 
-- Target Devices: 
-- Description: 
----------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity canvas is
    port (
        clk_i : in std_logic;
        write_enable_i : in std_logic;
        write_data_i : in std_logic_vector (0 to 79);
        write_address_i : in integer range 0 to 29;
        read_address_i : in integer range 0 to 29;
        read_data_o : out std_logic_vector (0 to 79)
    );
end canvas;

architecture Behavioral of canvas is
    type canvas_t is array (0 to 29) of std_logic_vector (0 to 79);
    signal canvas_data : canvas_t := (
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000011010101000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000001000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000001000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000001000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000001010100000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000001100000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000",
        "00000000000000000000000000000000000000000000000000000000000000000000000000000000"
    );
begin

    set : process( clk_i )
    begin
        if rising_edge( clk_i ) then
            if write_enable_i = '1' then
                canvas_data(write_address_i) <= write_data_i;
            end if ;
        end if ;
    end process ; -- set

    read_data_o <= canvas_data(read_address_i);

end Behavioral;